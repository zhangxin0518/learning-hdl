`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/06/18 20:54:36
// Design Name: 
// Module Name: tb_led_water
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_led_water(

    );                                           //Verilog��������ļ�û�������������

//----------------------------------------------------------------------------------------------------------------------------
reg clk;                                        //�����������ļ����������������һ���������������ģ��
reg datain;

//----------------------------------------------------------------------------------------------------------------------------
led_water   uut(                                //ʵ������������Ե��ļ���led_waterΪ������ģ�飬uutΪʵ����
    .clk(clk),                                  //���(���ұ�)Ϊ������ģ��Ľӿڣ��ұ�(�����ڱ���)Ϊ������ģ�鶨��ı���
    .datain(datain),
    .dataout(dataout)
);

//----------------------------------------------------------------------------------------------------------------------------
initial begin                                   //���д�������Ϊ������Լ��������д����
    clk <= 0;
    datain <= 0;
end

always #10 clk <= ~clk;
always #100 datain <= ~datain; 
    
endmodule






