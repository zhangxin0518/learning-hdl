// Verilog操作运算符
//---------------------------------------
1) 算术运算符(+,－,×，/,％) 
2) 赋值运算符(=,<=) 
3) 关系运算符(>,<,>=,<=,==,!=,===,!==) 
4) 逻辑运算符(&&,||,!) 
5) 条件运算符(?:) 
6) 位运算符(~,|,^,&,^~) 
7) 移位运算符(<<,>>) 
8) 拼接运算符({ })

// Verilog关键字
//----------------------------------------
always， and， assign，begin，buf，bufif0，
bufif1，case，casex，casez，cmos，deassign， 
default，defparam，disable，edge，else，end，
endcase，endmodule，endfunction，endprimitive, 
endspecify, endtable， endtask， event， for，
force， forever， fork， function，highz0，
highz1, if，initial, inout, input，integer，
join,large，macromodule，medium，module， nand，
negedge，nmos，nor，not，notif0，notifl, or, 
output, parameter, pmos, posedge, primitive, 
pull0, pull1, pullup, pulldown, rcmos, reg, 
releses, repeat, mmos, rpmos, rtran, rtranif0,
rtranif1,scalared,small，specify，specparam，
strength，strong0, strong1, supply0, supply1, 
table, task, time, tran, tranif0, tranif1, tri, 
tri0, tri1, triand, trior， trireg，vectored，
wait，wand，weak0，weak1，while， wire，wor, xnor，xor


